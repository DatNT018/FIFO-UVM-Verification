`ifndef FIFO_PARAM_PKG_SVH
`define FIFO_PARAM_PKG_SVH

package fifo_param_pkg;
	parameter FIFO_WIDTH = 4;
	parameter FIFO_DEPTH = 32;
	parameter FIFO_ADDR = 5;
endpackage

`endif
